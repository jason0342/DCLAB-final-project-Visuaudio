module IIRfilter(
	input i_clk,
	input i_rst
	// input i_data [31:0]fixpoint?
);