module DSP(
	input i_clk,
	input i_rst,
	input i_enable,
	input [15:0] i_data,
	output[15:0] o_data
);