module IIRfilter(
	input i_clk,
	input i_rst,
	input i_setparam,
	// input i_param [?:0]fixpoint?
	// input i_data [?:0]fixpoint?
);